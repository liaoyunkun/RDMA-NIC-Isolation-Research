module station_reader;
endmodule