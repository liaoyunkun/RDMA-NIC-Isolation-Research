`default_nettype none
`timescale 1ns/1ps

module slice_station;


endmodule